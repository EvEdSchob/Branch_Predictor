`timescale 1ns / 1ps

module BHT_1Bit(

    );
endmodule

`timescale 1ns / 1ps

module BHT_2Bit(

    );
endmodule